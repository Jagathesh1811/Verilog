module hs(input a, b, output d, br);
  assign d = a ^ b;
  assign br = ~a & b;
endmodule

